module CSAM(Z, X, Y);

        input logic [18:0] Y;
        input logic [18:0] X;
        output logic [37:0] Z;


        logic [18:0] P0;
        logic [18:0] carry1;
        logic [18:0] sum1;
        logic [18:0] P1;
        logic [18:0] carry2;
        logic [18:0] sum2;
        logic [18:0] P2;
        logic [18:0] carry3;
        logic [18:0] sum3;
        logic [18:0] P3;
        logic [18:0] carry4;
        logic [18:0] sum4;
        logic [18:0] P4;
        logic [18:0] carry5;
        logic [18:0] sum5;
        logic [18:0] P5;
        logic [18:0] carry6;
        logic [18:0] sum6;
        logic [18:0] P6;
        logic [18:0] carry7;
        logic [18:0] sum7;
        logic [18:0] P7;
        logic [18:0] carry8;
        logic [18:0] sum8;
        logic [18:0] P8;
        logic [18:0] carry9;
        logic [18:0] sum9;
        logic [18:0] P9;
        logic [18:0] carry10;
        logic [18:0] sum10;
        logic [18:0] P10;
        logic [18:0] carry11;
        logic [18:0] sum11;
        logic [18:0] P11;
        logic [18:0] carry12;
        logic [18:0] sum12;
        logic [18:0] P12;
        logic [18:0] carry13;
        logic [18:0] sum13;
        logic [18:0] P13;
        logic [18:0] carry14;
        logic [18:0] sum14;
        logic [18:0] P14;
        logic [18:0] carry15;
        logic [18:0] sum15;
        logic [18:0] P15;
        logic [18:0] carry16;
        logic [18:0] sum16;
        logic [18:0] P16;
        logic [18:0] carry17;
        logic [18:0] sum17;
        logic [18:0] P17;
        logic [18:0] carry18;
        logic [18:0] sum18;
        logic [18:0] P18;
        logic [18:0] carry19;
        logic [18:0] sum19;
        logic [36:0] carry20;


        // generate the partial products.
        partialProduct pp1(P0[18], X[18], Y[0]);
        partialProduct pp2(P0[17], X[17], Y[0]);
        partialProduct pp3(P0[16], X[16], Y[0]);
        partialProduct pp4(P0[15], X[15], Y[0]);
        partialProduct pp5(P0[14], X[14], Y[0]);
        partialProduct pp6(P0[13], X[13], Y[0]);
        partialProduct pp7(P0[12], X[12], Y[0]);
        partialProduct pp8(P0[11], X[11], Y[0]);
        partialProduct pp9(P0[10], X[10], Y[0]);
        partialProduct pp10(P0[9], X[9], Y[0]);
        partialProduct pp11(P0[8], X[8], Y[0]);
        partialProduct pp12(P0[7], X[7], Y[0]);
        partialProduct pp13(P0[6], X[6], Y[0]);
        partialProduct pp14(P0[5], X[5], Y[0]);
        partialProduct pp15(P0[4], X[4], Y[0]);
        partialProduct pp16(P0[3], X[3], Y[0]);
        partialProduct pp17(P0[2], X[2], Y[0]);
        partialProduct pp18(P0[1], X[1], Y[0]);
        partialProduct pp19(P0[0], X[0], Y[0]);
        partialProduct pp20(sum1[18], X[18], Y[1]);
        partialProduct pp21(P1[17], X[17], Y[1]);
        partialProduct pp22(P1[16], X[16], Y[1]);
        partialProduct pp23(P1[15], X[15], Y[1]);
        partialProduct pp24(P1[14], X[14], Y[1]);
        partialProduct pp25(P1[13], X[13], Y[1]);
        partialProduct pp26(P1[12], X[12], Y[1]);
        partialProduct pp27(P1[11], X[11], Y[1]);
        partialProduct pp28(P1[10], X[10], Y[1]);
        partialProduct pp29(P1[9], X[9], Y[1]);
        partialProduct pp30(P1[8], X[8], Y[1]);
        partialProduct pp31(P1[7], X[7], Y[1]);
        partialProduct pp32(P1[6], X[6], Y[1]);
        partialProduct pp33(P1[5], X[5], Y[1]);
        partialProduct pp34(P1[4], X[4], Y[1]);
        partialProduct pp35(P1[3], X[3], Y[1]);
        partialProduct pp36(P1[2], X[2], Y[1]);
        partialProduct pp37(P1[1], X[1], Y[1]);
        partialProduct pp38(P1[0], X[0], Y[1]);
        partialProduct pp39(sum2[18], X[18], Y[2]);
        partialProduct pp40(P2[17], X[17], Y[2]);
        partialProduct pp41(P2[16], X[16], Y[2]);
        partialProduct pp42(P2[15], X[15], Y[2]);
        partialProduct pp43(P2[14], X[14], Y[2]);
        partialProduct pp44(P2[13], X[13], Y[2]);
        partialProduct pp45(P2[12], X[12], Y[2]);
        partialProduct pp46(P2[11], X[11], Y[2]);
        partialProduct pp47(P2[10], X[10], Y[2]);
        partialProduct pp48(P2[9], X[9], Y[2]);
        partialProduct pp49(P2[8], X[8], Y[2]);
        partialProduct pp50(P2[7], X[7], Y[2]);
        partialProduct pp51(P2[6], X[6], Y[2]);
        partialProduct pp52(P2[5], X[5], Y[2]);
        partialProduct pp53(P2[4], X[4], Y[2]);
        partialProduct pp54(P2[3], X[3], Y[2]);
        partialProduct pp55(P2[2], X[2], Y[2]);
        partialProduct pp56(P2[1], X[1], Y[2]);
        partialProduct pp57(P2[0], X[0], Y[2]);
        partialProduct pp58(sum3[18], X[18], Y[3]);
        partialProduct pp59(P3[17], X[17], Y[3]);
        partialProduct pp60(P3[16], X[16], Y[3]);
        partialProduct pp61(P3[15], X[15], Y[3]);
        partialProduct pp62(P3[14], X[14], Y[3]);
        partialProduct pp63(P3[13], X[13], Y[3]);
        partialProduct pp64(P3[12], X[12], Y[3]);
        partialProduct pp65(P3[11], X[11], Y[3]);
        partialProduct pp66(P3[10], X[10], Y[3]);
        partialProduct pp67(P3[9], X[9], Y[3]);
        partialProduct pp68(P3[8], X[8], Y[3]);
        partialProduct pp69(P3[7], X[7], Y[3]);
        partialProduct pp70(P3[6], X[6], Y[3]);
        partialProduct pp71(P3[5], X[5], Y[3]);
        partialProduct pp72(P3[4], X[4], Y[3]);
        partialProduct pp73(P3[3], X[3], Y[3]);
        partialProduct pp74(P3[2], X[2], Y[3]);
        partialProduct pp75(P3[1], X[1], Y[3]);
        partialProduct pp76(P3[0], X[0], Y[3]);
        partialProduct pp77(sum4[18], X[18], Y[4]);
        partialProduct pp78(P4[17], X[17], Y[4]);
        partialProduct pp79(P4[16], X[16], Y[4]);
        partialProduct pp80(P4[15], X[15], Y[4]);
        partialProduct pp81(P4[14], X[14], Y[4]);
        partialProduct pp82(P4[13], X[13], Y[4]);
        partialProduct pp83(P4[12], X[12], Y[4]);
        partialProduct pp84(P4[11], X[11], Y[4]);
        partialProduct pp85(P4[10], X[10], Y[4]);
        partialProduct pp86(P4[9], X[9], Y[4]);
        partialProduct pp87(P4[8], X[8], Y[4]);
        partialProduct pp88(P4[7], X[7], Y[4]);
        partialProduct pp89(P4[6], X[6], Y[4]);
        partialProduct pp90(P4[5], X[5], Y[4]);
        partialProduct pp91(P4[4], X[4], Y[4]);
        partialProduct pp92(P4[3], X[3], Y[4]);
        partialProduct pp93(P4[2], X[2], Y[4]);
        partialProduct pp94(P4[1], X[1], Y[4]);
        partialProduct pp95(P4[0], X[0], Y[4]);
        partialProduct pp96(sum5[18], X[18], Y[5]);
        partialProduct pp97(P5[17], X[17], Y[5]);
        partialProduct pp98(P5[16], X[16], Y[5]);
        partialProduct pp99(P5[15], X[15], Y[5]);
        partialProduct pp100(P5[14], X[14], Y[5]);
        partialProduct pp101(P5[13], X[13], Y[5]);
        partialProduct pp102(P5[12], X[12], Y[5]);
        partialProduct pp103(P5[11], X[11], Y[5]);
        partialProduct pp104(P5[10], X[10], Y[5]);
        partialProduct pp105(P5[9], X[9], Y[5]);
        partialProduct pp106(P5[8], X[8], Y[5]);
        partialProduct pp107(P5[7], X[7], Y[5]);
        partialProduct pp108(P5[6], X[6], Y[5]);
        partialProduct pp109(P5[5], X[5], Y[5]);
        partialProduct pp110(P5[4], X[4], Y[5]);
        partialProduct pp111(P5[3], X[3], Y[5]);
        partialProduct pp112(P5[2], X[2], Y[5]);
        partialProduct pp113(P5[1], X[1], Y[5]);
        partialProduct pp114(P5[0], X[0], Y[5]);
        partialProduct pp115(sum6[18], X[18], Y[6]);
        partialProduct pp116(P6[17], X[17], Y[6]);
        partialProduct pp117(P6[16], X[16], Y[6]);
        partialProduct pp118(P6[15], X[15], Y[6]);
        partialProduct pp119(P6[14], X[14], Y[6]);
        partialProduct pp120(P6[13], X[13], Y[6]);
        partialProduct pp121(P6[12], X[12], Y[6]);
        partialProduct pp122(P6[11], X[11], Y[6]);
        partialProduct pp123(P6[10], X[10], Y[6]);
        partialProduct pp124(P6[9], X[9], Y[6]);
        partialProduct pp125(P6[8], X[8], Y[6]);
        partialProduct pp126(P6[7], X[7], Y[6]);
        partialProduct pp127(P6[6], X[6], Y[6]);
        partialProduct pp128(P6[5], X[5], Y[6]);
        partialProduct pp129(P6[4], X[4], Y[6]);
        partialProduct pp130(P6[3], X[3], Y[6]);
        partialProduct pp131(P6[2], X[2], Y[6]);
        partialProduct pp132(P6[1], X[1], Y[6]);
        partialProduct pp133(P6[0], X[0], Y[6]);
        partialProduct pp134(sum7[18], X[18], Y[7]);
        partialProduct pp135(P7[17], X[17], Y[7]);
        partialProduct pp136(P7[16], X[16], Y[7]);
        partialProduct pp137(P7[15], X[15], Y[7]);
        partialProduct pp138(P7[14], X[14], Y[7]);
        partialProduct pp139(P7[13], X[13], Y[7]);
        partialProduct pp140(P7[12], X[12], Y[7]);
        partialProduct pp141(P7[11], X[11], Y[7]);
        partialProduct pp142(P7[10], X[10], Y[7]);
        partialProduct pp143(P7[9], X[9], Y[7]);
        partialProduct pp144(P7[8], X[8], Y[7]);
        partialProduct pp145(P7[7], X[7], Y[7]);
        partialProduct pp146(P7[6], X[6], Y[7]);
        partialProduct pp147(P7[5], X[5], Y[7]);
        partialProduct pp148(P7[4], X[4], Y[7]);
        partialProduct pp149(P7[3], X[3], Y[7]);
        partialProduct pp150(P7[2], X[2], Y[7]);
        partialProduct pp151(P7[1], X[1], Y[7]);
        partialProduct pp152(P7[0], X[0], Y[7]);
        partialProduct pp153(sum8[18], X[18], Y[8]);
        partialProduct pp154(P8[17], X[17], Y[8]);
        partialProduct pp155(P8[16], X[16], Y[8]);
        partialProduct pp156(P8[15], X[15], Y[8]);
        partialProduct pp157(P8[14], X[14], Y[8]);
        partialProduct pp158(P8[13], X[13], Y[8]);
        partialProduct pp159(P8[12], X[12], Y[8]);
        partialProduct pp160(P8[11], X[11], Y[8]);
        partialProduct pp161(P8[10], X[10], Y[8]);
        partialProduct pp162(P8[9], X[9], Y[8]);
        partialProduct pp163(P8[8], X[8], Y[8]);
        partialProduct pp164(P8[7], X[7], Y[8]);
        partialProduct pp165(P8[6], X[6], Y[8]);
        partialProduct pp166(P8[5], X[5], Y[8]);
        partialProduct pp167(P8[4], X[4], Y[8]);
        partialProduct pp168(P8[3], X[3], Y[8]);
        partialProduct pp169(P8[2], X[2], Y[8]);
        partialProduct pp170(P8[1], X[1], Y[8]);
        partialProduct pp171(P8[0], X[0], Y[8]);
        partialProduct pp172(sum9[18], X[18], Y[9]);
        partialProduct pp173(P9[17], X[17], Y[9]);
        partialProduct pp174(P9[16], X[16], Y[9]);
        partialProduct pp175(P9[15], X[15], Y[9]);
        partialProduct pp176(P9[14], X[14], Y[9]);
        partialProduct pp177(P9[13], X[13], Y[9]);
        partialProduct pp178(P9[12], X[12], Y[9]);
        partialProduct pp179(P9[11], X[11], Y[9]);
        partialProduct pp180(P9[10], X[10], Y[9]);
        partialProduct pp181(P9[9], X[9], Y[9]);
        partialProduct pp182(P9[8], X[8], Y[9]);
        partialProduct pp183(P9[7], X[7], Y[9]);
        partialProduct pp184(P9[6], X[6], Y[9]);
        partialProduct pp185(P9[5], X[5], Y[9]);
        partialProduct pp186(P9[4], X[4], Y[9]);
        partialProduct pp187(P9[3], X[3], Y[9]);
        partialProduct pp188(P9[2], X[2], Y[9]);
        partialProduct pp189(P9[1], X[1], Y[9]);
        partialProduct pp190(P9[0], X[0], Y[9]);
        partialProduct pp191(sum10[18], X[18], Y[10]);
        partialProduct pp192(P10[17], X[17], Y[10]);
        partialProduct pp193(P10[16], X[16], Y[10]);
        partialProduct pp194(P10[15], X[15], Y[10]);
        partialProduct pp195(P10[14], X[14], Y[10]);
        partialProduct pp196(P10[13], X[13], Y[10]);
        partialProduct pp197(P10[12], X[12], Y[10]);
        partialProduct pp198(P10[11], X[11], Y[10]);
        partialProduct pp199(P10[10], X[10], Y[10]);
        partialProduct pp200(P10[9], X[9], Y[10]);
        partialProduct pp201(P10[8], X[8], Y[10]);
        partialProduct pp202(P10[7], X[7], Y[10]);
        partialProduct pp203(P10[6], X[6], Y[10]);
        partialProduct pp204(P10[5], X[5], Y[10]);
        partialProduct pp205(P10[4], X[4], Y[10]);
        partialProduct pp206(P10[3], X[3], Y[10]);
        partialProduct pp207(P10[2], X[2], Y[10]);
        partialProduct pp208(P10[1], X[1], Y[10]);
        partialProduct pp209(P10[0], X[0], Y[10]);
        partialProduct pp210(sum11[18], X[18], Y[11]);
        partialProduct pp211(P11[17], X[17], Y[11]);
        partialProduct pp212(P11[16], X[16], Y[11]);
        partialProduct pp213(P11[15], X[15], Y[11]);
        partialProduct pp214(P11[14], X[14], Y[11]);
        partialProduct pp215(P11[13], X[13], Y[11]);
        partialProduct pp216(P11[12], X[12], Y[11]);
        partialProduct pp217(P11[11], X[11], Y[11]);
        partialProduct pp218(P11[10], X[10], Y[11]);
        partialProduct pp219(P11[9], X[9], Y[11]);
        partialProduct pp220(P11[8], X[8], Y[11]);
        partialProduct pp221(P11[7], X[7], Y[11]);
        partialProduct pp222(P11[6], X[6], Y[11]);
        partialProduct pp223(P11[5], X[5], Y[11]);
        partialProduct pp224(P11[4], X[4], Y[11]);
        partialProduct pp225(P11[3], X[3], Y[11]);
        partialProduct pp226(P11[2], X[2], Y[11]);
        partialProduct pp227(P11[1], X[1], Y[11]);
        partialProduct pp228(P11[0], X[0], Y[11]);
        partialProduct pp229(sum12[18], X[18], Y[12]);
        partialProduct pp230(P12[17], X[17], Y[12]);
        partialProduct pp231(P12[16], X[16], Y[12]);
        partialProduct pp232(P12[15], X[15], Y[12]);
        partialProduct pp233(P12[14], X[14], Y[12]);
        partialProduct pp234(P12[13], X[13], Y[12]);
        partialProduct pp235(P12[12], X[12], Y[12]);
        partialProduct pp236(P12[11], X[11], Y[12]);
        partialProduct pp237(P12[10], X[10], Y[12]);
        partialProduct pp238(P12[9], X[9], Y[12]);
        partialProduct pp239(P12[8], X[8], Y[12]);
        partialProduct pp240(P12[7], X[7], Y[12]);
        partialProduct pp241(P12[6], X[6], Y[12]);
        partialProduct pp242(P12[5], X[5], Y[12]);
        partialProduct pp243(P12[4], X[4], Y[12]);
        partialProduct pp244(P12[3], X[3], Y[12]);
        partialProduct pp245(P12[2], X[2], Y[12]);
        partialProduct pp246(P12[1], X[1], Y[12]);
        partialProduct pp247(P12[0], X[0], Y[12]);
        partialProduct pp248(sum13[18], X[18], Y[13]);
        partialProduct pp249(P13[17], X[17], Y[13]);
        partialProduct pp250(P13[16], X[16], Y[13]);
        partialProduct pp251(P13[15], X[15], Y[13]);
        partialProduct pp252(P13[14], X[14], Y[13]);
        partialProduct pp253(P13[13], X[13], Y[13]);
        partialProduct pp254(P13[12], X[12], Y[13]);
        partialProduct pp255(P13[11], X[11], Y[13]);
        partialProduct pp256(P13[10], X[10], Y[13]);
        partialProduct pp257(P13[9], X[9], Y[13]);
        partialProduct pp258(P13[8], X[8], Y[13]);
        partialProduct pp259(P13[7], X[7], Y[13]);
        partialProduct pp260(P13[6], X[6], Y[13]);
        partialProduct pp261(P13[5], X[5], Y[13]);
        partialProduct pp262(P13[4], X[4], Y[13]);
        partialProduct pp263(P13[3], X[3], Y[13]);
        partialProduct pp264(P13[2], X[2], Y[13]);
        partialProduct pp265(P13[1], X[1], Y[13]);
        partialProduct pp266(P13[0], X[0], Y[13]);
        partialProduct pp267(sum14[18], X[18], Y[14]);
        partialProduct pp268(P14[17], X[17], Y[14]);
        partialProduct pp269(P14[16], X[16], Y[14]);
        partialProduct pp270(P14[15], X[15], Y[14]);
        partialProduct pp271(P14[14], X[14], Y[14]);
        partialProduct pp272(P14[13], X[13], Y[14]);
        partialProduct pp273(P14[12], X[12], Y[14]);
        partialProduct pp274(P14[11], X[11], Y[14]);
        partialProduct pp275(P14[10], X[10], Y[14]);
        partialProduct pp276(P14[9], X[9], Y[14]);
        partialProduct pp277(P14[8], X[8], Y[14]);
        partialProduct pp278(P14[7], X[7], Y[14]);
        partialProduct pp279(P14[6], X[6], Y[14]);
        partialProduct pp280(P14[5], X[5], Y[14]);
        partialProduct pp281(P14[4], X[4], Y[14]);
        partialProduct pp282(P14[3], X[3], Y[14]);
        partialProduct pp283(P14[2], X[2], Y[14]);
        partialProduct pp284(P14[1], X[1], Y[14]);
        partialProduct pp285(P14[0], X[0], Y[14]);
        partialProduct pp286(sum15[18], X[18], Y[15]);
        partialProduct pp287(P15[17], X[17], Y[15]);
        partialProduct pp288(P15[16], X[16], Y[15]);
        partialProduct pp289(P15[15], X[15], Y[15]);
        partialProduct pp290(P15[14], X[14], Y[15]);
        partialProduct pp291(P15[13], X[13], Y[15]);
        partialProduct pp292(P15[12], X[12], Y[15]);
        partialProduct pp293(P15[11], X[11], Y[15]);
        partialProduct pp294(P15[10], X[10], Y[15]);
        partialProduct pp295(P15[9], X[9], Y[15]);
        partialProduct pp296(P15[8], X[8], Y[15]);
        partialProduct pp297(P15[7], X[7], Y[15]);
        partialProduct pp298(P15[6], X[6], Y[15]);
        partialProduct pp299(P15[5], X[5], Y[15]);
        partialProduct pp300(P15[4], X[4], Y[15]);
        partialProduct pp301(P15[3], X[3], Y[15]);
        partialProduct pp302(P15[2], X[2], Y[15]);
        partialProduct pp303(P15[1], X[1], Y[15]);
        partialProduct pp304(P15[0], X[0], Y[15]);
        partialProduct pp305(sum16[18], X[18], Y[16]);
        partialProduct pp306(P16[17], X[17], Y[16]);
        partialProduct pp307(P16[16], X[16], Y[16]);
        partialProduct pp308(P16[15], X[15], Y[16]);
        partialProduct pp309(P16[14], X[14], Y[16]);
        partialProduct pp310(P16[13], X[13], Y[16]);
        partialProduct pp311(P16[12], X[12], Y[16]);
        partialProduct pp312(P16[11], X[11], Y[16]);
        partialProduct pp313(P16[10], X[10], Y[16]);
        partialProduct pp314(P16[9], X[9], Y[16]);
        partialProduct pp315(P16[8], X[8], Y[16]);
        partialProduct pp316(P16[7], X[7], Y[16]);
        partialProduct pp317(P16[6], X[6], Y[16]);
        partialProduct pp318(P16[5], X[5], Y[16]);
        partialProduct pp319(P16[4], X[4], Y[16]);
        partialProduct pp320(P16[3], X[3], Y[16]);
        partialProduct pp321(P16[2], X[2], Y[16]);
        partialProduct pp322(P16[1], X[1], Y[16]);
        partialProduct pp323(P16[0], X[0], Y[16]);
        partialProduct pp324(sum17[18], X[18], Y[17]);
        partialProduct pp325(P17[17], X[17], Y[17]);
        partialProduct pp326(P17[16], X[16], Y[17]);
        partialProduct pp327(P17[15], X[15], Y[17]);
        partialProduct pp328(P17[14], X[14], Y[17]);
        partialProduct pp329(P17[13], X[13], Y[17]);
        partialProduct pp330(P17[12], X[12], Y[17]);
        partialProduct pp331(P17[11], X[11], Y[17]);
        partialProduct pp332(P17[10], X[10], Y[17]);
        partialProduct pp333(P17[9], X[9], Y[17]);
        partialProduct pp334(P17[8], X[8], Y[17]);
        partialProduct pp335(P17[7], X[7], Y[17]);
        partialProduct pp336(P17[6], X[6], Y[17]);
        partialProduct pp337(P17[5], X[5], Y[17]);
        partialProduct pp338(P17[4], X[4], Y[17]);
        partialProduct pp339(P17[3], X[3], Y[17]);
        partialProduct pp340(P17[2], X[2], Y[17]);
        partialProduct pp341(P17[1], X[1], Y[17]);
        partialProduct pp342(P17[0], X[0], Y[17]);
        partialProduct pp343(sum18[18], X[18], Y[18]);
        partialProduct pp344(P18[17], X[17], Y[18]);
        partialProduct pp345(P18[16], X[16], Y[18]);
        partialProduct pp346(P18[15], X[15], Y[18]);
        partialProduct pp347(P18[14], X[14], Y[18]);
        partialProduct pp348(P18[13], X[13], Y[18]);
        partialProduct pp349(P18[12], X[12], Y[18]);
        partialProduct pp350(P18[11], X[11], Y[18]);
        partialProduct pp351(P18[10], X[10], Y[18]);
        partialProduct pp352(P18[9], X[9], Y[18]);
        partialProduct pp353(P18[8], X[8], Y[18]);
        partialProduct pp354(P18[7], X[7], Y[18]);
        partialProduct pp355(P18[6], X[6], Y[18]);
        partialProduct pp356(P18[5], X[5], Y[18]);
        partialProduct pp357(P18[4], X[4], Y[18]);
        partialProduct pp358(P18[3], X[3], Y[18]);
        partialProduct pp359(P18[2], X[2], Y[18]);
        partialProduct pp360(P18[1], X[1], Y[18]);
        partialProduct pp361(P18[0], X[0], Y[18]);

        // Array Reduction
        half_adder  HA1(carry1[17],sum1[17],P1[17],P0[18]);
        half_adder  HA2(carry1[16],sum1[16],P1[16],P0[17]);
        half_adder  HA3(carry1[15],sum1[15],P1[15],P0[16]);
        half_adder  HA4(carry1[14],sum1[14],P1[14],P0[15]);
        half_adder  HA5(carry1[13],sum1[13],P1[13],P0[14]);
        half_adder  HA6(carry1[12],sum1[12],P1[12],P0[13]);
        half_adder  HA7(carry1[11],sum1[11],P1[11],P0[12]);
        half_adder  HA8(carry1[10],sum1[10],P1[10],P0[11]);
        half_adder  HA9(carry1[9],sum1[9],P1[9],P0[10]);
        half_adder  HA10(carry1[8],sum1[8],P1[8],P0[9]);
        half_adder  HA11(carry1[7],sum1[7],P1[7],P0[8]);
        half_adder  HA12(carry1[6],sum1[6],P1[6],P0[7]);
        half_adder  HA13(carry1[5],sum1[5],P1[5],P0[6]);
        half_adder  HA14(carry1[4],sum1[4],P1[4],P0[5]);
        half_adder  HA15(carry1[3],sum1[3],P1[3],P0[4]);
        half_adder  HA16(carry1[2],sum1[2],P1[2],P0[3]);
        half_adder  HA17(carry1[1],sum1[1],P1[1],P0[2]);
        half_adder  HA18(carry1[0],sum1[0],P1[0],P0[1]);
        full_adder  FA1(carry2[17],sum2[17],P2[17],sum1[18],carry1[17]);
        full_adder  FA2(carry2[16],sum2[16],P2[16],sum1[17],carry1[16]);
        full_adder  FA3(carry2[15],sum2[15],P2[15],sum1[16],carry1[15]);
        full_adder  FA4(carry2[14],sum2[14],P2[14],sum1[15],carry1[14]);
        full_adder  FA5(carry2[13],sum2[13],P2[13],sum1[14],carry1[13]);
        full_adder  FA6(carry2[12],sum2[12],P2[12],sum1[13],carry1[12]);
        full_adder  FA7(carry2[11],sum2[11],P2[11],sum1[12],carry1[11]);
        full_adder  FA8(carry2[10],sum2[10],P2[10],sum1[11],carry1[10]);
        full_adder  FA9(carry2[9],sum2[9],P2[9],sum1[10],carry1[9]);
        full_adder  FA10(carry2[8],sum2[8],P2[8],sum1[9],carry1[8]);
        full_adder  FA11(carry2[7],sum2[7],P2[7],sum1[8],carry1[7]);
        full_adder  FA12(carry2[6],sum2[6],P2[6],sum1[7],carry1[6]);
        full_adder  FA13(carry2[5],sum2[5],P2[5],sum1[6],carry1[5]);
        full_adder  FA14(carry2[4],sum2[4],P2[4],sum1[5],carry1[4]);
        full_adder  FA15(carry2[3],sum2[3],P2[3],sum1[4],carry1[3]);
        full_adder  FA16(carry2[2],sum2[2],P2[2],sum1[3],carry1[2]);
        full_adder  FA17(carry2[1],sum2[1],P2[1],sum1[2],carry1[1]);
        full_adder  FA18(carry2[0],sum2[0],P2[0],sum1[1],carry1[0]);
        full_adder  FA19(carry3[17],sum3[17],P3[17],sum2[18],carry2[17]);
        full_adder  FA20(carry3[16],sum3[16],P3[16],sum2[17],carry2[16]);
        full_adder  FA21(carry3[15],sum3[15],P3[15],sum2[16],carry2[15]);
        full_adder  FA22(carry3[14],sum3[14],P3[14],sum2[15],carry2[14]);
        full_adder  FA23(carry3[13],sum3[13],P3[13],sum2[14],carry2[13]);
        full_adder  FA24(carry3[12],sum3[12],P3[12],sum2[13],carry2[12]);
        full_adder  FA25(carry3[11],sum3[11],P3[11],sum2[12],carry2[11]);
        full_adder  FA26(carry3[10],sum3[10],P3[10],sum2[11],carry2[10]);
        full_adder  FA27(carry3[9],sum3[9],P3[9],sum2[10],carry2[9]);
        full_adder  FA28(carry3[8],sum3[8],P3[8],sum2[9],carry2[8]);
        full_adder  FA29(carry3[7],sum3[7],P3[7],sum2[8],carry2[7]);
        full_adder  FA30(carry3[6],sum3[6],P3[6],sum2[7],carry2[6]);
        full_adder  FA31(carry3[5],sum3[5],P3[5],sum2[6],carry2[5]);
        full_adder  FA32(carry3[4],sum3[4],P3[4],sum2[5],carry2[4]);
        full_adder  FA33(carry3[3],sum3[3],P3[3],sum2[4],carry2[3]);
        full_adder  FA34(carry3[2],sum3[2],P3[2],sum2[3],carry2[2]);
        full_adder  FA35(carry3[1],sum3[1],P3[1],sum2[2],carry2[1]);
        full_adder  FA36(carry3[0],sum3[0],P3[0],sum2[1],carry2[0]);
        full_adder  FA37(carry4[17],sum4[17],P4[17],sum3[18],carry3[17]);
        full_adder  FA38(carry4[16],sum4[16],P4[16],sum3[17],carry3[16]);
        full_adder  FA39(carry4[15],sum4[15],P4[15],sum3[16],carry3[15]);
        full_adder  FA40(carry4[14],sum4[14],P4[14],sum3[15],carry3[14]);
        full_adder  FA41(carry4[13],sum4[13],P4[13],sum3[14],carry3[13]);
        full_adder  FA42(carry4[12],sum4[12],P4[12],sum3[13],carry3[12]);
        full_adder  FA43(carry4[11],sum4[11],P4[11],sum3[12],carry3[11]);
        full_adder  FA44(carry4[10],sum4[10],P4[10],sum3[11],carry3[10]);
        full_adder  FA45(carry4[9],sum4[9],P4[9],sum3[10],carry3[9]);
        full_adder  FA46(carry4[8],sum4[8],P4[8],sum3[9],carry3[8]);
        full_adder  FA47(carry4[7],sum4[7],P4[7],sum3[8],carry3[7]);
        full_adder  FA48(carry4[6],sum4[6],P4[6],sum3[7],carry3[6]);
        full_adder  FA49(carry4[5],sum4[5],P4[5],sum3[6],carry3[5]);
        full_adder  FA50(carry4[4],sum4[4],P4[4],sum3[5],carry3[4]);
        full_adder  FA51(carry4[3],sum4[3],P4[3],sum3[4],carry3[3]);
        full_adder  FA52(carry4[2],sum4[2],P4[2],sum3[3],carry3[2]);
        full_adder  FA53(carry4[1],sum4[1],P4[1],sum3[2],carry3[1]);
        full_adder  FA54(carry4[0],sum4[0],P4[0],sum3[1],carry3[0]);
        full_adder  FA55(carry5[17],sum5[17],P5[17],sum4[18],carry4[17]);
        full_adder  FA56(carry5[16],sum5[16],P5[16],sum4[17],carry4[16]);
        full_adder  FA57(carry5[15],sum5[15],P5[15],sum4[16],carry4[15]);
        full_adder  FA58(carry5[14],sum5[14],P5[14],sum4[15],carry4[14]);
        full_adder  FA59(carry5[13],sum5[13],P5[13],sum4[14],carry4[13]);
        full_adder  FA60(carry5[12],sum5[12],P5[12],sum4[13],carry4[12]);
        full_adder  FA61(carry5[11],sum5[11],P5[11],sum4[12],carry4[11]);
        full_adder  FA62(carry5[10],sum5[10],P5[10],sum4[11],carry4[10]);
        full_adder  FA63(carry5[9],sum5[9],P5[9],sum4[10],carry4[9]);
        full_adder  FA64(carry5[8],sum5[8],P5[8],sum4[9],carry4[8]);
        full_adder  FA65(carry5[7],sum5[7],P5[7],sum4[8],carry4[7]);
        full_adder  FA66(carry5[6],sum5[6],P5[6],sum4[7],carry4[6]);
        full_adder  FA67(carry5[5],sum5[5],P5[5],sum4[6],carry4[5]);
        full_adder  FA68(carry5[4],sum5[4],P5[4],sum4[5],carry4[4]);
        full_adder  FA69(carry5[3],sum5[3],P5[3],sum4[4],carry4[3]);
        full_adder  FA70(carry5[2],sum5[2],P5[2],sum4[3],carry4[2]);
        full_adder  FA71(carry5[1],sum5[1],P5[1],sum4[2],carry4[1]);
        full_adder  FA72(carry5[0],sum5[0],P5[0],sum4[1],carry4[0]);
        full_adder  FA73(carry6[17],sum6[17],P6[17],sum5[18],carry5[17]);
        full_adder  FA74(carry6[16],sum6[16],P6[16],sum5[17],carry5[16]);
        full_adder  FA75(carry6[15],sum6[15],P6[15],sum5[16],carry5[15]);
        full_adder  FA76(carry6[14],sum6[14],P6[14],sum5[15],carry5[14]);
        full_adder  FA77(carry6[13],sum6[13],P6[13],sum5[14],carry5[13]);
        full_adder  FA78(carry6[12],sum6[12],P6[12],sum5[13],carry5[12]);
        full_adder  FA79(carry6[11],sum6[11],P6[11],sum5[12],carry5[11]);
        full_adder  FA80(carry6[10],sum6[10],P6[10],sum5[11],carry5[10]);
        full_adder  FA81(carry6[9],sum6[9],P6[9],sum5[10],carry5[9]);
        full_adder  FA82(carry6[8],sum6[8],P6[8],sum5[9],carry5[8]);
        full_adder  FA83(carry6[7],sum6[7],P6[7],sum5[8],carry5[7]);
        full_adder  FA84(carry6[6],sum6[6],P6[6],sum5[7],carry5[6]);
        full_adder  FA85(carry6[5],sum6[5],P6[5],sum5[6],carry5[5]);
        full_adder  FA86(carry6[4],sum6[4],P6[4],sum5[5],carry5[4]);
        full_adder  FA87(carry6[3],sum6[3],P6[3],sum5[4],carry5[3]);
        full_adder  FA88(carry6[2],sum6[2],P6[2],sum5[3],carry5[2]);
        full_adder  FA89(carry6[1],sum6[1],P6[1],sum5[2],carry5[1]);
        full_adder  FA90(carry6[0],sum6[0],P6[0],sum5[1],carry5[0]);
        full_adder  FA91(carry7[17],sum7[17],P7[17],sum6[18],carry6[17]);
        full_adder  FA92(carry7[16],sum7[16],P7[16],sum6[17],carry6[16]);
        full_adder  FA93(carry7[15],sum7[15],P7[15],sum6[16],carry6[15]);
        full_adder  FA94(carry7[14],sum7[14],P7[14],sum6[15],carry6[14]);
        full_adder  FA95(carry7[13],sum7[13],P7[13],sum6[14],carry6[13]);
        full_adder  FA96(carry7[12],sum7[12],P7[12],sum6[13],carry6[12]);
        full_adder  FA97(carry7[11],sum7[11],P7[11],sum6[12],carry6[11]);
        full_adder  FA98(carry7[10],sum7[10],P7[10],sum6[11],carry6[10]);
        full_adder  FA99(carry7[9],sum7[9],P7[9],sum6[10],carry6[9]);
        full_adder  FA100(carry7[8],sum7[8],P7[8],sum6[9],carry6[8]);
        full_adder  FA101(carry7[7],sum7[7],P7[7],sum6[8],carry6[7]);
        full_adder  FA102(carry7[6],sum7[6],P7[6],sum6[7],carry6[6]);
        full_adder  FA103(carry7[5],sum7[5],P7[5],sum6[6],carry6[5]);
        full_adder  FA104(carry7[4],sum7[4],P7[4],sum6[5],carry6[4]);
        full_adder  FA105(carry7[3],sum7[3],P7[3],sum6[4],carry6[3]);
        full_adder  FA106(carry7[2],sum7[2],P7[2],sum6[3],carry6[2]);
        full_adder  FA107(carry7[1],sum7[1],P7[1],sum6[2],carry6[1]);
        full_adder  FA108(carry7[0],sum7[0],P7[0],sum6[1],carry6[0]);
        full_adder  FA109(carry8[17],sum8[17],P8[17],sum7[18],carry7[17]);
        full_adder  FA110(carry8[16],sum8[16],P8[16],sum7[17],carry7[16]);
        full_adder  FA111(carry8[15],sum8[15],P8[15],sum7[16],carry7[15]);
        full_adder  FA112(carry8[14],sum8[14],P8[14],sum7[15],carry7[14]);
        full_adder  FA113(carry8[13],sum8[13],P8[13],sum7[14],carry7[13]);
        full_adder  FA114(carry8[12],sum8[12],P8[12],sum7[13],carry7[12]);
        full_adder  FA115(carry8[11],sum8[11],P8[11],sum7[12],carry7[11]);
        full_adder  FA116(carry8[10],sum8[10],P8[10],sum7[11],carry7[10]);
        full_adder  FA117(carry8[9],sum8[9],P8[9],sum7[10],carry7[9]);
        full_adder  FA118(carry8[8],sum8[8],P8[8],sum7[9],carry7[8]);
        full_adder  FA119(carry8[7],sum8[7],P8[7],sum7[8],carry7[7]);
        full_adder  FA120(carry8[6],sum8[6],P8[6],sum7[7],carry7[6]);
        full_adder  FA121(carry8[5],sum8[5],P8[5],sum7[6],carry7[5]);
        full_adder  FA122(carry8[4],sum8[4],P8[4],sum7[5],carry7[4]);
        full_adder  FA123(carry8[3],sum8[3],P8[3],sum7[4],carry7[3]);
        full_adder  FA124(carry8[2],sum8[2],P8[2],sum7[3],carry7[2]);
        full_adder  FA125(carry8[1],sum8[1],P8[1],sum7[2],carry7[1]);
        full_adder  FA126(carry8[0],sum8[0],P8[0],sum7[1],carry7[0]);
        full_adder  FA127(carry9[17],sum9[17],P9[17],sum8[18],carry8[17]);
        full_adder  FA128(carry9[16],sum9[16],P9[16],sum8[17],carry8[16]);
        full_adder  FA129(carry9[15],sum9[15],P9[15],sum8[16],carry8[15]);
        full_adder  FA130(carry9[14],sum9[14],P9[14],sum8[15],carry8[14]);
        full_adder  FA131(carry9[13],sum9[13],P9[13],sum8[14],carry8[13]);
        full_adder  FA132(carry9[12],sum9[12],P9[12],sum8[13],carry8[12]);
        full_adder  FA133(carry9[11],sum9[11],P9[11],sum8[12],carry8[11]);
        full_adder  FA134(carry9[10],sum9[10],P9[10],sum8[11],carry8[10]);
        full_adder  FA135(carry9[9],sum9[9],P9[9],sum8[10],carry8[9]);
        full_adder  FA136(carry9[8],sum9[8],P9[8],sum8[9],carry8[8]);
        full_adder  FA137(carry9[7],sum9[7],P9[7],sum8[8],carry8[7]);
        full_adder  FA138(carry9[6],sum9[6],P9[6],sum8[7],carry8[6]);
        full_adder  FA139(carry9[5],sum9[5],P9[5],sum8[6],carry8[5]);
        full_adder  FA140(carry9[4],sum9[4],P9[4],sum8[5],carry8[4]);
        full_adder  FA141(carry9[3],sum9[3],P9[3],sum8[4],carry8[3]);
        full_adder  FA142(carry9[2],sum9[2],P9[2],sum8[3],carry8[2]);
        full_adder  FA143(carry9[1],sum9[1],P9[1],sum8[2],carry8[1]);
        full_adder  FA144(carry9[0],sum9[0],P9[0],sum8[1],carry8[0]);
        full_adder  FA145(carry10[17],sum10[17],P10[17],sum9[18],carry9[17]);
        full_adder  FA146(carry10[16],sum10[16],P10[16],sum9[17],carry9[16]);
        full_adder  FA147(carry10[15],sum10[15],P10[15],sum9[16],carry9[15]);
        full_adder  FA148(carry10[14],sum10[14],P10[14],sum9[15],carry9[14]);
        full_adder  FA149(carry10[13],sum10[13],P10[13],sum9[14],carry9[13]);
        full_adder  FA150(carry10[12],sum10[12],P10[12],sum9[13],carry9[12]);
        full_adder  FA151(carry10[11],sum10[11],P10[11],sum9[12],carry9[11]);
        full_adder  FA152(carry10[10],sum10[10],P10[10],sum9[11],carry9[10]);
        full_adder  FA153(carry10[9],sum10[9],P10[9],sum9[10],carry9[9]);
        full_adder  FA154(carry10[8],sum10[8],P10[8],sum9[9],carry9[8]);
        full_adder  FA155(carry10[7],sum10[7],P10[7],sum9[8],carry9[7]);
        full_adder  FA156(carry10[6],sum10[6],P10[6],sum9[7],carry9[6]);
        full_adder  FA157(carry10[5],sum10[5],P10[5],sum9[6],carry9[5]);
        full_adder  FA158(carry10[4],sum10[4],P10[4],sum9[5],carry9[4]);
        full_adder  FA159(carry10[3],sum10[3],P10[3],sum9[4],carry9[3]);
        full_adder  FA160(carry10[2],sum10[2],P10[2],sum9[3],carry9[2]);
        full_adder  FA161(carry10[1],sum10[1],P10[1],sum9[2],carry9[1]);
        full_adder  FA162(carry10[0],sum10[0],P10[0],sum9[1],carry9[0]);
        full_adder  FA163(carry11[17],sum11[17],P11[17],sum10[18],carry10[17]);
        full_adder  FA164(carry11[16],sum11[16],P11[16],sum10[17],carry10[16]);
        full_adder  FA165(carry11[15],sum11[15],P11[15],sum10[16],carry10[15]);
        full_adder  FA166(carry11[14],sum11[14],P11[14],sum10[15],carry10[14]);
        full_adder  FA167(carry11[13],sum11[13],P11[13],sum10[14],carry10[13]);
        full_adder  FA168(carry11[12],sum11[12],P11[12],sum10[13],carry10[12]);
        full_adder  FA169(carry11[11],sum11[11],P11[11],sum10[12],carry10[11]);
        full_adder  FA170(carry11[10],sum11[10],P11[10],sum10[11],carry10[10]);
        full_adder  FA171(carry11[9],sum11[9],P11[9],sum10[10],carry10[9]);
        full_adder  FA172(carry11[8],sum11[8],P11[8],sum10[9],carry10[8]);
        full_adder  FA173(carry11[7],sum11[7],P11[7],sum10[8],carry10[7]);
        full_adder  FA174(carry11[6],sum11[6],P11[6],sum10[7],carry10[6]);
        full_adder  FA175(carry11[5],sum11[5],P11[5],sum10[6],carry10[5]);
        full_adder  FA176(carry11[4],sum11[4],P11[4],sum10[5],carry10[4]);
        full_adder  FA177(carry11[3],sum11[3],P11[3],sum10[4],carry10[3]);
        full_adder  FA178(carry11[2],sum11[2],P11[2],sum10[3],carry10[2]);
        full_adder  FA179(carry11[1],sum11[1],P11[1],sum10[2],carry10[1]);
        full_adder  FA180(carry11[0],sum11[0],P11[0],sum10[1],carry10[0]);
        full_adder  FA181(carry12[17],sum12[17],P12[17],sum11[18],carry11[17]);
        full_adder  FA182(carry12[16],sum12[16],P12[16],sum11[17],carry11[16]);
        full_adder  FA183(carry12[15],sum12[15],P12[15],sum11[16],carry11[15]);
        full_adder  FA184(carry12[14],sum12[14],P12[14],sum11[15],carry11[14]);
        full_adder  FA185(carry12[13],sum12[13],P12[13],sum11[14],carry11[13]);
        full_adder  FA186(carry12[12],sum12[12],P12[12],sum11[13],carry11[12]);
        full_adder  FA187(carry12[11],sum12[11],P12[11],sum11[12],carry11[11]);
        full_adder  FA188(carry12[10],sum12[10],P12[10],sum11[11],carry11[10]);
        full_adder  FA189(carry12[9],sum12[9],P12[9],sum11[10],carry11[9]);
        full_adder  FA190(carry12[8],sum12[8],P12[8],sum11[9],carry11[8]);
        full_adder  FA191(carry12[7],sum12[7],P12[7],sum11[8],carry11[7]);
        full_adder  FA192(carry12[6],sum12[6],P12[6],sum11[7],carry11[6]);
        full_adder  FA193(carry12[5],sum12[5],P12[5],sum11[6],carry11[5]);
        full_adder  FA194(carry12[4],sum12[4],P12[4],sum11[5],carry11[4]);
        full_adder  FA195(carry12[3],sum12[3],P12[3],sum11[4],carry11[3]);
        full_adder  FA196(carry12[2],sum12[2],P12[2],sum11[3],carry11[2]);
        full_adder  FA197(carry12[1],sum12[1],P12[1],sum11[2],carry11[1]);
        full_adder  FA198(carry12[0],sum12[0],P12[0],sum11[1],carry11[0]);
        full_adder  FA199(carry13[17],sum13[17],P13[17],sum12[18],carry12[17]);
        full_adder  FA200(carry13[16],sum13[16],P13[16],sum12[17],carry12[16]);
        full_adder  FA201(carry13[15],sum13[15],P13[15],sum12[16],carry12[15]);
        full_adder  FA202(carry13[14],sum13[14],P13[14],sum12[15],carry12[14]);
        full_adder  FA203(carry13[13],sum13[13],P13[13],sum12[14],carry12[13]);
        full_adder  FA204(carry13[12],sum13[12],P13[12],sum12[13],carry12[12]);
        full_adder  FA205(carry13[11],sum13[11],P13[11],sum12[12],carry12[11]);
        full_adder  FA206(carry13[10],sum13[10],P13[10],sum12[11],carry12[10]);
        full_adder  FA207(carry13[9],sum13[9],P13[9],sum12[10],carry12[9]);
        full_adder  FA208(carry13[8],sum13[8],P13[8],sum12[9],carry12[8]);
        full_adder  FA209(carry13[7],sum13[7],P13[7],sum12[8],carry12[7]);
        full_adder  FA210(carry13[6],sum13[6],P13[6],sum12[7],carry12[6]);
        full_adder  FA211(carry13[5],sum13[5],P13[5],sum12[6],carry12[5]);
        full_adder  FA212(carry13[4],sum13[4],P13[4],sum12[5],carry12[4]);
        full_adder  FA213(carry13[3],sum13[3],P13[3],sum12[4],carry12[3]);
        full_adder  FA214(carry13[2],sum13[2],P13[2],sum12[3],carry12[2]);
        full_adder  FA215(carry13[1],sum13[1],P13[1],sum12[2],carry12[1]);
        full_adder  FA216(carry13[0],sum13[0],P13[0],sum12[1],carry12[0]);
        full_adder  FA217(carry14[17],sum14[17],P14[17],sum13[18],carry13[17]);
        full_adder  FA218(carry14[16],sum14[16],P14[16],sum13[17],carry13[16]);
        full_adder  FA219(carry14[15],sum14[15],P14[15],sum13[16],carry13[15]);
        full_adder  FA220(carry14[14],sum14[14],P14[14],sum13[15],carry13[14]);
        full_adder  FA221(carry14[13],sum14[13],P14[13],sum13[14],carry13[13]);
        full_adder  FA222(carry14[12],sum14[12],P14[12],sum13[13],carry13[12]);
        full_adder  FA223(carry14[11],sum14[11],P14[11],sum13[12],carry13[11]);
        full_adder  FA224(carry14[10],sum14[10],P14[10],sum13[11],carry13[10]);
        full_adder  FA225(carry14[9],sum14[9],P14[9],sum13[10],carry13[9]);
        full_adder  FA226(carry14[8],sum14[8],P14[8],sum13[9],carry13[8]);
        full_adder  FA227(carry14[7],sum14[7],P14[7],sum13[8],carry13[7]);
        full_adder  FA228(carry14[6],sum14[6],P14[6],sum13[7],carry13[6]);
        full_adder  FA229(carry14[5],sum14[5],P14[5],sum13[6],carry13[5]);
        full_adder  FA230(carry14[4],sum14[4],P14[4],sum13[5],carry13[4]);
        full_adder  FA231(carry14[3],sum14[3],P14[3],sum13[4],carry13[3]);
        full_adder  FA232(carry14[2],sum14[2],P14[2],sum13[3],carry13[2]);
        full_adder  FA233(carry14[1],sum14[1],P14[1],sum13[2],carry13[1]);
        full_adder  FA234(carry14[0],sum14[0],P14[0],sum13[1],carry13[0]);
        full_adder  FA235(carry15[17],sum15[17],P15[17],sum14[18],carry14[17]);
        full_adder  FA236(carry15[16],sum15[16],P15[16],sum14[17],carry14[16]);
        full_adder  FA237(carry15[15],sum15[15],P15[15],sum14[16],carry14[15]);
        full_adder  FA238(carry15[14],sum15[14],P15[14],sum14[15],carry14[14]);
        full_adder  FA239(carry15[13],sum15[13],P15[13],sum14[14],carry14[13]);
        full_adder  FA240(carry15[12],sum15[12],P15[12],sum14[13],carry14[12]);
        full_adder  FA241(carry15[11],sum15[11],P15[11],sum14[12],carry14[11]);
        full_adder  FA242(carry15[10],sum15[10],P15[10],sum14[11],carry14[10]);
        full_adder  FA243(carry15[9],sum15[9],P15[9],sum14[10],carry14[9]);
        full_adder  FA244(carry15[8],sum15[8],P15[8],sum14[9],carry14[8]);
        full_adder  FA245(carry15[7],sum15[7],P15[7],sum14[8],carry14[7]);
        full_adder  FA246(carry15[6],sum15[6],P15[6],sum14[7],carry14[6]);
        full_adder  FA247(carry15[5],sum15[5],P15[5],sum14[6],carry14[5]);
        full_adder  FA248(carry15[4],sum15[4],P15[4],sum14[5],carry14[4]);
        full_adder  FA249(carry15[3],sum15[3],P15[3],sum14[4],carry14[3]);
        full_adder  FA250(carry15[2],sum15[2],P15[2],sum14[3],carry14[2]);
        full_adder  FA251(carry15[1],sum15[1],P15[1],sum14[2],carry14[1]);
        full_adder  FA252(carry15[0],sum15[0],P15[0],sum14[1],carry14[0]);
        full_adder  FA253(carry16[17],sum16[17],P16[17],sum15[18],carry15[17]);
        full_adder  FA254(carry16[16],sum16[16],P16[16],sum15[17],carry15[16]);
        full_adder  FA255(carry16[15],sum16[15],P16[15],sum15[16],carry15[15]);
        full_adder  FA256(carry16[14],sum16[14],P16[14],sum15[15],carry15[14]);
        full_adder  FA257(carry16[13],sum16[13],P16[13],sum15[14],carry15[13]);
        full_adder  FA258(carry16[12],sum16[12],P16[12],sum15[13],carry15[12]);
        full_adder  FA259(carry16[11],sum16[11],P16[11],sum15[12],carry15[11]);
        full_adder  FA260(carry16[10],sum16[10],P16[10],sum15[11],carry15[10]);
        full_adder  FA261(carry16[9],sum16[9],P16[9],sum15[10],carry15[9]);
        full_adder  FA262(carry16[8],sum16[8],P16[8],sum15[9],carry15[8]);
        full_adder  FA263(carry16[7],sum16[7],P16[7],sum15[8],carry15[7]);
        full_adder  FA264(carry16[6],sum16[6],P16[6],sum15[7],carry15[6]);
        full_adder  FA265(carry16[5],sum16[5],P16[5],sum15[6],carry15[5]);
        full_adder  FA266(carry16[4],sum16[4],P16[4],sum15[5],carry15[4]);
        full_adder  FA267(carry16[3],sum16[3],P16[3],sum15[4],carry15[3]);
        full_adder  FA268(carry16[2],sum16[2],P16[2],sum15[3],carry15[2]);
        full_adder  FA269(carry16[1],sum16[1],P16[1],sum15[2],carry15[1]);
        full_adder  FA270(carry16[0],sum16[0],P16[0],sum15[1],carry15[0]);
        full_adder  FA271(carry17[17],sum17[17],P17[17],sum16[18],carry16[17]);
        full_adder  FA272(carry17[16],sum17[16],P17[16],sum16[17],carry16[16]);
        full_adder  FA273(carry17[15],sum17[15],P17[15],sum16[16],carry16[15]);
        full_adder  FA274(carry17[14],sum17[14],P17[14],sum16[15],carry16[14]);
        full_adder  FA275(carry17[13],sum17[13],P17[13],sum16[14],carry16[13]);
        full_adder  FA276(carry17[12],sum17[12],P17[12],sum16[13],carry16[12]);
        full_adder  FA277(carry17[11],sum17[11],P17[11],sum16[12],carry16[11]);
        full_adder  FA278(carry17[10],sum17[10],P17[10],sum16[11],carry16[10]);
        full_adder  FA279(carry17[9],sum17[9],P17[9],sum16[10],carry16[9]);
        full_adder  FA280(carry17[8],sum17[8],P17[8],sum16[9],carry16[8]);
        full_adder  FA281(carry17[7],sum17[7],P17[7],sum16[8],carry16[7]);
        full_adder  FA282(carry17[6],sum17[6],P17[6],sum16[7],carry16[6]);
        full_adder  FA283(carry17[5],sum17[5],P17[5],sum16[6],carry16[5]);
        full_adder  FA284(carry17[4],sum17[4],P17[4],sum16[5],carry16[4]);
        full_adder  FA285(carry17[3],sum17[3],P17[3],sum16[4],carry16[3]);
        full_adder  FA286(carry17[2],sum17[2],P17[2],sum16[3],carry16[2]);
        full_adder  FA287(carry17[1],sum17[1],P17[1],sum16[2],carry16[1]);
        full_adder  FA288(carry17[0],sum17[0],P17[0],sum16[1],carry16[0]);
        full_adder  FA289(carry18[17],sum18[17],P18[17],sum17[18],carry17[17]);
        full_adder  FA290(carry18[16],sum18[16],P18[16],sum17[17],carry17[16]);
        full_adder  FA291(carry18[15],sum18[15],P18[15],sum17[16],carry17[15]);
        full_adder  FA292(carry18[14],sum18[14],P18[14],sum17[15],carry17[14]);
        full_adder  FA293(carry18[13],sum18[13],P18[13],sum17[14],carry17[13]);
        full_adder  FA294(carry18[12],sum18[12],P18[12],sum17[13],carry17[12]);
        full_adder  FA295(carry18[11],sum18[11],P18[11],sum17[12],carry17[11]);
        full_adder  FA296(carry18[10],sum18[10],P18[10],sum17[11],carry17[10]);
        full_adder  FA297(carry18[9],sum18[9],P18[9],sum17[10],carry17[9]);
        full_adder  FA298(carry18[8],sum18[8],P18[8],sum17[9],carry17[8]);
        full_adder  FA299(carry18[7],sum18[7],P18[7],sum17[8],carry17[7]);
        full_adder  FA300(carry18[6],sum18[6],P18[6],sum17[7],carry17[6]);
        full_adder  FA301(carry18[5],sum18[5],P18[5],sum17[6],carry17[5]);
        full_adder  FA302(carry18[4],sum18[4],P18[4],sum17[5],carry17[4]);
        full_adder  FA303(carry18[3],sum18[3],P18[3],sum17[4],carry17[3]);
        full_adder  FA304(carry18[2],sum18[2],P18[2],sum17[3],carry17[2]);
        full_adder  FA305(carry18[1],sum18[1],P18[1],sum17[2],carry17[1]);
        full_adder  FA306(carry18[0],sum18[0],P18[0],sum17[1],carry17[0]);

        // Generate lower product bits YBITS
        buf b1(Z[0], P0[0]);
        assign Z[1] = sum1[0];
        assign Z[2] = sum2[0];
        assign Z[3] = sum3[0];
        assign Z[4] = sum4[0];
        assign Z[5] = sum5[0];
        assign Z[6] = sum6[0];
        assign Z[7] = sum7[0];
        assign Z[8] = sum8[0];
        assign Z[9] = sum9[0];
        assign Z[10] = sum10[0];
        assign Z[11] = sum11[0];
        assign Z[12] = sum12[0];
        assign Z[13] = sum13[0];
        assign Z[14] = sum14[0];
        assign Z[15] = sum15[0];
        assign Z[16] = sum16[0];
        assign Z[17] = sum17[0];
        assign Z[18] = sum18[0];

        // Final Carry Propagate Addition
        half_adder CPA1(carry19[0],Z[19],carry18[0],sum18[1]);
        full_adder CPA2(carry19[1],Z[20],carry18[1],carry19[0],sum18[2]);
        full_adder CPA3(carry19[2],Z[21],carry18[2],carry19[1],sum18[3]);
        full_adder CPA4(carry19[3],Z[22],carry18[3],carry19[2],sum18[4]);
        full_adder CPA5(carry19[4],Z[23],carry18[4],carry19[3],sum18[5]);
        full_adder CPA6(carry19[5],Z[24],carry18[5],carry19[4],sum18[6]);
        full_adder CPA7(carry19[6],Z[25],carry18[6],carry19[5],sum18[7]);
        full_adder CPA8(carry19[7],Z[26],carry18[7],carry19[6],sum18[8]);
        full_adder CPA9(carry19[8],Z[27],carry18[8],carry19[7],sum18[9]);
        full_adder CPA10(carry19[9],Z[28],carry18[9],carry19[8],sum18[10]);
        full_adder CPA11(carry19[10],Z[29],carry18[10],carry19[9],sum18[11]);
        full_adder CPA12(carry19[11],Z[30],carry18[11],carry19[10],sum18[12]);
        full_adder CPA13(carry19[12],Z[31],carry18[12],carry19[11],sum18[13]);
        full_adder CPA14(carry19[13],Z[32],carry18[13],carry19[12],sum18[14]);
        full_adder CPA15(carry19[14],Z[33],carry18[14],carry19[13],sum18[15]);
        full_adder CPA16(carry19[15],Z[34],carry18[15],carry19[14],sum18[16]);
        full_adder CPA17(carry19[16],Z[35],carry18[16],carry19[15],sum18[17]);
        full_adder CPA18(Z[37],Z[36],carry18[17],carry19[16],sum18[18]);

endmodule
