module RNE(input logic[31:0] big,
            output logic [15:0] rounded);

endmodule
