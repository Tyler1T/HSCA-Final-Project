module and3 (input logic a, b, c,
                output logic out);

endmodule // and3
