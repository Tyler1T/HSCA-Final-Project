module flipper (input logic a,
            output logic notA);

    assign notA = ~a;

endmodule // not
