module mux4by16(input  logic [15:0]     d0, d1, d2, d3,
                input  logic [1:0]      S,
                output logic [15:0]     Y);

    mux4 m0 (Y[0], d0[0], d1[0], d2[0], d3[0], S);
    mux4 m1 (Y[1], d0[1], d1[1], d2[1], d3[1], S);
    mux4 m2 (Y[2], d0[2], d1[2], d2[2], d3[2], S);
    mux4 m3 (Y[3], d0[3], d1[3], d2[3], d3[3], S);
    mux4 m4 (Y[4], d0[4], d1[4], d2[4], d3[4], S);
    mux4 m5 (Y[5], d0[5], d1[5], d2[5], d3[5], S);
    mux4 m6 (Y[6], d0[6], d1[6], d2[6], d3[6], S);
    mux4 m7 (Y[7], d0[7], d1[7], d2[7], d3[7], S);
    mux4 m8 (Y[8], d0[8], d1[8], d2[8], d3[8], S);
    mux4 m9 (Y[9], d0[9], d1[9], d2[9], d3[9], S);
    mux4 m10 (Y[10], d0[10], d1[10], d2[10], d3[10], S);
    mux4 m11 (Y[11], d0[11], d1[11], d2[11], d3[11], S);
    mux4 m12 (Y[12], d0[12], d1[12], d2[12], d3[12], S);
    mux4 m13 (Y[13], d0[13], d1[13], d2[13], d3[13], S);
    mux4 m14 (Y[14], d0[14], d1[14], d2[14], d3[14], S);
    mux4 m15 (Y[15], d0[15], d1[15], d2[15], d3[15], S);


endmodule // mux41
